module _4zm16Selector (clk, rst, \�_____ , A3, A2, A1, A0, \0 , \1 , \2 , \3 , \4 , \5 , \6 , \7 , \8 , \9 , A, B, C, D, E, F);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [0:0] \�_____ ;
  input  wire [0:0] A3;
  input  wire [0:0] A2;
  input  wire [0:0] A1;
  input  wire [0:0] A0;
  output  wire [0:0] \0 ;
  output  wire [0:0] \1 ;
  output  wire [0:0] \2 ;
  output  wire [0:0] \3 ;
  output  wire [0:0] \4 ;
  output  wire [0:0] \5 ;
  output  wire [0:0] \6 ;
  output  wire [0:0] \7 ;
  output  wire [0:0] \8 ;
  output  wire [0:0] \9 ;
  output  wire [0:0] A;
  output  wire [0:0] B;
  output  wire [0:0] C;
  output  wire [0:0] D;
  output  wire [0:0] E;
  output  wire [0:0] F;

  TC_Decoder3 # (.UUID(64'd2564989398389830754 ^ UUID)) Decoder3_0 (.dis(wire_17), .sel0(wire_6), .sel1(wire_9), .sel2(wire_1), .out0(wire_11), .out1(wire_12), .out2(wire_20), .out3(wire_3), .out4(wire_10), .out5(wire_23), .out6(wire_21), .out7(wire_15));
  TC_Decoder3 # (.UUID(64'd2298840035739462038 ^ UUID)) Decoder3_1 (.dis(wire_5), .sel0(wire_6), .sel1(wire_9), .sel2(wire_1), .out0(wire_22), .out1(wire_8), .out2(wire_13), .out3(wire_2), .out4(wire_19), .out5(wire_7), .out6(wire_14), .out7(wire_18));
  TC_Or # (.UUID(64'd3175078524024449064 ^ UUID), .BIT_WIDTH(64'd1)) Or_2 (.in0(wire_4), .in1(wire_0), .out(wire_5));
  TC_Not # (.UUID(64'd2061859652610692002 ^ UUID), .BIT_WIDTH(64'd1)) Not_3 (.in(wire_4), .out(wire_16));
  TC_Or # (.UUID(64'd1447438233748301576 ^ UUID), .BIT_WIDTH(64'd1)) Or_4 (.in0(wire_16), .in1(wire_0), .out(wire_17));
  TC_Constant # (.UUID(64'd4553024698181830824 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_5 (.out());
  TC_Constant # (.UUID(64'd2064339905802656346 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_6 (.out());
  TC_Constant # (.UUID(64'd2735987545437809334 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_7 (.out());
  TC_Constant # (.UUID(64'd879239978781978394 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_8 (.out());
  TC_Constant # (.UUID(64'd3030286631431832873 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_9 (.out());
  TC_Constant # (.UUID(64'd3261601882157773873 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_10 (.out());
  TC_Constant # (.UUID(64'd2854776969465089937 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_11 (.out());
  TC_Constant # (.UUID(64'd871924067805957400 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_12 (.out());
  TC_Constant # (.UUID(64'd3260889488327193501 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_13 (.out());
  TC_Constant # (.UUID(64'd486451695951613651 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_14 (.out());
  TC_Constant # (.UUID(64'd2551029110425735131 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_15 (.out());
  TC_Constant # (.UUID(64'd3824417624477149852 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_16 (.out());
  TC_Constant # (.UUID(64'd4219020160871176370 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_17 (.out());
  TC_Constant # (.UUID(64'd1080587990143207529 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_18 (.out());
  TC_Constant # (.UUID(64'd2188918196940788858 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_19 (.out());
  TC_Constant # (.UUID(64'd4449410397033879695 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_20 (.out());
  TC_Constant # (.UUID(64'd683406866284922864 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_21 (.out());
  TC_Constant # (.UUID(64'd1092000694853377679 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_22 (.out());
  TC_Constant # (.UUID(64'd654324742496264292 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_23 (.out());
  TC_Constant # (.UUID(64'd3131037719329940983 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_24 (.out());
  TC_Constant # (.UUID(64'd3704327759118139311 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_25 (.out());
  TC_Constant # (.UUID(64'd2786119359103655322 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_26 (.out());
  TC_Constant # (.UUID(64'd4547717834180229615 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_27 (.out());
  TC_Constant # (.UUID(64'd1360817414555130003 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_28 (.out());
  TC_Constant # (.UUID(64'd378917427681715807 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_29 (.out());

  wire [0:0] wire_0;
  assign wire_0 = \�_____ ;
  wire [0:0] wire_1;
  assign wire_1 = A2;
  wire [0:0] wire_2;
  assign \3  = wire_2;
  wire [0:0] wire_3;
  assign B = wire_3;
  wire [0:0] wire_4;
  assign wire_4 = A3;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  assign wire_6 = A0;
  wire [0:0] wire_7;
  assign \5  = wire_7;
  wire [0:0] wire_8;
  assign \1  = wire_8;
  wire [0:0] wire_9;
  assign wire_9 = A1;
  wire [0:0] wire_10;
  assign C = wire_10;
  wire [0:0] wire_11;
  assign \8  = wire_11;
  wire [0:0] wire_12;
  assign \9  = wire_12;
  wire [0:0] wire_13;
  assign \2  = wire_13;
  wire [0:0] wire_14;
  assign \6  = wire_14;
  wire [0:0] wire_15;
  assign F = wire_15;
  wire [0:0] wire_16;
  wire [0:0] wire_17;
  wire [0:0] wire_18;
  assign \7  = wire_18;
  wire [0:0] wire_19;
  assign \4  = wire_19;
  wire [0:0] wire_20;
  assign A = wire_20;
  wire [0:0] wire_21;
  assign E = wire_21;
  wire [0:0] wire_22;
  assign \0  = wire_22;
  wire [0:0] wire_23;
  assign D = wire_23;

endmodule
