module HfcloudzmLEG (clk, rst, arch_output_enable, arch_output_value, arch_input_enable, arch_input_value);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  output  wire [0:0] arch_output_enable;
  output  wire [7:0] arch_output_value;
  output  wire [0:0] arch_input_enable;
  input  wire [7:0] arch_input_value;

  TC_IOSwitch # (.UUID(64'd4389593845 ^ UUID), .BIT_WIDTH(64'd8)) LevelOutputArch_0 (.in(wire_31), .en(wire_87), .out(arch_output_value));
  TC_Constant # (.UUID(64'd646894894600596568 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h6)) Constant8_1 (.out(wire_38));
  TC_Constant # (.UUID(64'd1561870452110776218 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h7)) Constant8_2 (.out(wire_20));
  TC_Equal # (.UUID(64'd1203356891022513320 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_3 (.in0(wire_38), .in1(wire_13[7:0]), .out(wire_16));
  TC_Equal # (.UUID(64'd1442812294779791168 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_4 (.in0(wire_38), .in1(wire_6[7:0]), .out(wire_61));
  TC_Equal # (.UUID(64'd2015717940966090344 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_5 (.in0(wire_20), .in1(wire_13[7:0]), .out(wire_4));
  TC_Equal # (.UUID(64'd406854493208215620 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_6 (.in0(wire_20), .in1(wire_6[7:0]), .out(wire_56));
  TC_Or # (.UUID(64'd231608398890168832 ^ UUID), .BIT_WIDTH(64'd1)) Or_7 (.in0(wire_4), .in1(wire_56), .out(wire_57));
  TC_Constant # (.UUID(64'd1146358017678501326 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h7)) Constant8_8 (.out(wire_58));
  TC_Equal # (.UUID(64'd3858704228872944971 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_9 (.in0(wire_3), .in1(wire_58), .out(wire_87));
  TC_Constant # (.UUID(64'd2452001502727780469 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h6)) Constant8_10 (.out(wire_74));
  TC_Mux # (.UUID(64'd3901832152078863778 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_11 (.sel(wire_84), .in0(wire_71), .in1(wire_13[7:0]), .out(wire_1));
  TC_Mux # (.UUID(64'd3459404181720251683 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_12 (.sel(wire_90), .in0(wire_76), .in1(wire_6[7:0]), .out(wire_27));
  TC_Splitter8 # (.UUID(64'd4039262554454177485 ^ UUID)) Splitter8_13 (.in(wire_10[7:0]), .out0(wire_11), .out1(wire_64), .out2(wire_48), .out3(), .out4(wire_82), .out5(wire_88), .out6(), .out7());
  TC_Maker8 # (.UUID(64'd490613999964465760 ^ UUID)) Maker8_14 (.in0(wire_11), .in1(wire_64), .in2(wire_48), .in3(1'd0), .in4(1'd0), .in5(1'd0), .in6(1'd0), .in7(1'd0), .out(wire_85));
  TC_And # (.UUID(64'd444835506320179650 ^ UUID), .BIT_WIDTH(64'd1)) And_15 (.in0(wire_67), .in1(wire_21), .out(wire_45));
  TC_Switch # (.UUID(64'd1690711706184722343 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_16 (.en(wire_18), .in(wire_5[7:0]), .out(wire_3));
  TC_Mux # (.UUID(64'd2250560463839008046 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_17 (.sel(wire_45), .in0(wire_31), .in1(wire_36), .out(wire_22));
  TC_Splitter8 # (.UUID(64'd3595891711551887685 ^ UUID)) Splitter8_18 (.in(wire_10[7:0]), .out0(wire_32), .out1(), .out2(), .out3(), .out4(wire_49), .out5(wire_54), .out6(), .out7());
  TC_Mux # (.UUID(64'd989258781171139647 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_19 (.sel(wire_50), .in0(wire_24), .in1(wire_46[7:0]), .out(wire_31));
  TC_And # (.UUID(64'd2963477707908923054 ^ UUID), .BIT_WIDTH(64'd1)) And_20 (.in0(wire_23), .in1(wire_2), .out(wire_50));
  TC_Not # (.UUID(64'd2945859350466821452 ^ UUID), .BIT_WIDTH(64'd1)) Not_21 (.in(wire_32), .out(wire_23));
  TC_And # (.UUID(64'd1041448334109548536 ^ UUID), .BIT_WIDTH(64'd1)) And_22 (.in0(wire_32), .in1(wire_2), .out(wire_53));
  TC_Or # (.UUID(64'd3444792903697950215 ^ UUID), .BIT_WIDTH(64'd1)) Or_23 (.in0(wire_50), .in1(wire_53), .out(wire_35));
  TC_Switch # (.UUID(64'd353561922716362211 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_24 (.en(wire_35), .in(wire_27), .out(wire_73));
  TC_Not # (.UUID(64'd1085057617843046386 ^ UUID), .BIT_WIDTH(64'd1)) Not_25 (.in(wire_53), .out(wire_40));
  TC_Not # (.UUID(64'd1510224717874120443 ^ UUID), .BIT_WIDTH(64'd1)) Not_26 (.in(wire_67), .out(wire_18));
  TC_Not # (.UUID(64'd3779063054668046542 ^ UUID), .BIT_WIDTH(64'd1)) Not_27 (.in(wire_54), .out(wire_72));
  TC_And # (.UUID(64'd146387254429518226 ^ UUID), .BIT_WIDTH(64'd1)) And_28 (.in0(wire_49), .in1(wire_72), .out(wire_2));
  TC_Not # (.UUID(64'd3566342795601416862 ^ UUID), .BIT_WIDTH(64'd1)) Not_29 (.in(wire_82), .out(wire_77));
  TC_And # (.UUID(64'd149690425414889478 ^ UUID), .BIT_WIDTH(64'd1)) And_30 (.in0(wire_77), .in1(wire_88), .out(wire_67));
  TC_Not # (.UUID(64'd3137639030705816530 ^ UUID), .BIT_WIDTH(64'd1)) Not_31 (.in(wire_14), .out(wire_42));
  TC_Not # (.UUID(64'd3035321497610409034 ^ UUID), .BIT_WIDTH(64'd1)) Not_32 (.in(wire_62), .out(wire_75));
  TC_And # (.UUID(64'd1540713049143640502 ^ UUID), .BIT_WIDTH(64'd1)) And_33 (.in0(wire_42), .in1(wire_75), .out(wire_52));
  TC_Mux # (.UUID(64'd2502500774298529496 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_34 (.sel(wire_52), .in0(wire_68), .in1(wire_30), .out(wire_24));
  TC_And # (.UUID(64'd1778810683900461498 ^ UUID), .BIT_WIDTH(64'd1)) And_35 (.in0(wire_37), .in1(wire_44), .out(wire_0));
  TC_Not # (.UUID(64'd412372632254406258 ^ UUID), .BIT_WIDTH(64'd1)) Not_36 (.in(wire_25), .out(wire_60));
  TC_And # (.UUID(64'd756821310729295725 ^ UUID), .BIT_WIDTH(64'd1)) And_37 (.in0(wire_60), .in1(wire_0), .out(wire_29));
  TC_And # (.UUID(64'd2524197232253226030 ^ UUID), .BIT_WIDTH(64'd1)) And_38 (.in0(wire_25), .in1(wire_0), .out(wire_47));
  TC_Add # (.UUID(64'd1658730676323503364 ^ UUID), .BIT_WIDTH(64'd8)) Add8_39 (.in0(wire_1), .in1(wire_81), .ci(1'd0), .out(wire_12), .co());
  TC_Constant # (.UUID(64'd1887338667276813868 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h4)) Constant8_40 (.out(wire_81));
  TC_Mux # (.UUID(64'd1016629334141804913 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_41 (.sel(wire_26), .in0(wire_1), .in1(wire_12), .out(wire_91));
  TC_Switch # (.UUID(64'd438959385 ^ UUID), .BIT_WIDTH(64'd8)) LevelInputArch_42 (.en(wire_57), .in(arch_input_value), .out(wire_70));
  TC_Counter # (.UUID(64'd812697445171396358 ^ UUID), .BIT_WIDTH(64'd8), .count(8'd4)) Counter8_43 (.clk(clk), .rst(rst), .save(wire_17), .in(wire_28), .out(wire_8));
  TC_Equal # (.UUID(64'd827106679222120445 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_44 (.in0(wire_74), .in1(wire_3), .out(wire_15));
  TC_Maker8 # (.UUID(64'd3738195046192671420 ^ UUID)) Maker8_45 (.in0(wire_51), .in1(wire_59), .in2(wire_43), .in3(wire_89), .in4(1'd0), .in5(1'd0), .in6(1'd0), .in7(1'd0), .out(wire_66));
  TC_Splitter8 # (.UUID(64'd1057503288219103610 ^ UUID)) Splitter8_46 (.in(wire_10[7:0]), .out0(wire_51), .out1(wire_59), .out2(wire_43), .out3(wire_89), .out4(wire_14), .out5(wire_62), .out6(wire_90), .out7(wire_84));
  TC_Splitter8 # (.UUID(64'd4508525212144124302 ^ UUID)) Splitter8_47 (.in(wire_10[7:0]), .out0(wire_25), .out1(wire_26), .out2(wire_19), .out3(), .out4(wire_37), .out5(wire_44), .out6(), .out7());
  TC_Ram # (.UUID(64'd4545406246428990035 ^ UUID), .WORD_WIDTH(64'd8), .WORD_COUNT(64'd256)) Ram_48 (.clk(clk), .rst(rst), .load(wire_50), .save(wire_53), .address({{24{1'b0}}, wire_73 }), .in0({{56{1'b0}}, wire_1 }), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_46), .out1(), .out2(), .out3());
  TC_Program # (.UUID(64'd3369947834646235778 ^ UUID), .WORD_WIDTH(64'd8), .DEFAULT_FILE_NAME("Program_2EC475B36BAF8A82.w8.bin"), .ARG_SIG("Program_2EC475B36BAF8A82=%s")) Program_49 (.clk(clk), .rst(rst), .address({{8{1'b0}}, wire_8 }), .out0(wire_10), .out1(wire_13), .out2(wire_6), .out3(wire_5));
  TC_And # (.UUID(64'd1594903537683014851 ^ UUID), .BIT_WIDTH(64'd1)) And_50 (.in0(wire_0), .in1(wire_7), .out(wire_9));
  TC_Or # (.UUID(64'd1489425258395036641 ^ UUID), .BIT_WIDTH(64'd1)) Or_51 (.in0(wire_19), .in1(wire_26), .out(wire_7));
  TC_Mux # (.UUID(64'd1960894067275396396 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_52 (.sel(wire_9), .in0(wire_22), .in1(wire_36), .out(wire_28));
  TC_Or3 # (.UUID(64'd2500749203645481152 ^ UUID), .BIT_WIDTH(64'd1)) Or3_53 (.in0(wire_15), .in1(wire_9), .in2(wire_45), .out(wire_17));
  TC_And # (.UUID(64'd2949321221645705801 ^ UUID), .BIT_WIDTH(64'd1)) And_54 (.in0(wire_0), .in1(wire_19), .out(wire_41));
  TC_Mux # (.UUID(64'd1242918659469910056 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_55 (.sel(wire_41), .in0(wire_5[7:0]), .in1(wire_33), .out(wire_36));
  TC_And3 # (.UUID(64'd2450443017567893698 ^ UUID), .BIT_WIDTH(64'd1)) And3_56 (.in0(wire_18), .in1(wire_34), .in2(wire_40), .out(wire_83));
  TC_Not # (.UUID(64'd3044943248572491271 ^ UUID), .BIT_WIDTH(64'd1)) Not_57 (.in(wire_41), .out(wire_34));
  TC_And # (.UUID(64'd610971993186129457 ^ UUID), .BIT_WIDTH(64'd1)) And_58 (.in0(wire_0), .in1(wire_26), .out(wire_65));
  TC_Not # (.UUID(64'd3494257868534462216 ^ UUID), .BIT_WIDTH(64'd1)) Not_59 (.in(wire_65), .out(wire_86));
  LEG_ALU # (.UUID(64'd1708942249613249991 ^ UUID)) LEG_ALU_60 (.clk(clk), .rst(rst), .OPCODE(wire_66), .OP1(wire_1), .OP2(wire_27), .Output(wire_30));
  LEG_COND # (.UUID(64'd392033239601748503 ^ UUID)) LEG_COND_61 (.clk(clk), .rst(rst), .OP1(wire_1), .OP2(wire_27), .OP(wire_85), .Output(wire_21));
  _3WayzmMUXzm8b # (.UUID(64'd3620365979226132878 ^ UUID)) _3WayzmMUXzm8b_62 (.clk(clk), .rst(rst), .In0(wire_69), .In1_1(wire_8), .In2_1(wire_70), .In1_2(wire_61), .In2_2(wire_56), .Out(wire_76));
  _3WayzmMUXzm8b # (.UUID(64'd1990550809129563582 ^ UUID)) _3WayzmMUXzm8b_63 (.clk(clk), .rst(rst), .In0(wire_39), .In1_1(wire_8), .In2_1(wire_70), .In1_2(wire_16), .In2_2(wire_4), .Out(wire_71));
  Stackzm8b # (.UUID(64'd4423945735032464992 ^ UUID)) Stackzm8b_64 (.clk(clk), .rst(rst), .POP(wire_47), .PUSH(wire_29), .VALUE(wire_91), .OUTPUT(wire_68), .Top(wire_33));
  RegisterFiles4x4zm8bzmEX # (.UUID(64'd483272188785477457 ^ UUID)) RegisterFiles4x4zm8bzmEX_65 (.clk(clk), .rst(rst), .R_ADDR2(wire_6[7:0]), .R_ADDR1(wire_13[7:0]), .\input (wire_31), .W(wire_80), .W_ADDR(wire_3), .READ_2(wire_69), .READ_1(wire_39));
  TC_Not # (.UUID(64'd3126466636152228092 ^ UUID), .BIT_WIDTH(64'd1)) Not_66 (.in(wire_25), .out(wire_78));
  TC_Not # (.UUID(64'd3809689304776512617 ^ UUID), .BIT_WIDTH(64'd1)) Not_67 (.in(wire_26), .out(wire_79));
  TC_And3 # (.UUID(64'd4610694646076225075 ^ UUID), .BIT_WIDTH(64'd1)) And3_68 (.in0(wire_0), .in1(wire_79), .in2(wire_78), .out(wire_55));
  TC_And3 # (.UUID(64'd177528929341615137 ^ UUID), .BIT_WIDTH(64'd1)) And3_69 (.in0(wire_83), .in1(wire_63), .in2(wire_86), .out(wire_80));
  TC_Not # (.UUID(64'd4157073821873738745 ^ UUID), .BIT_WIDTH(64'd1)) Not_70 (.in(wire_55), .out(wire_63));

  wire [0:0] wire_0;
  wire [7:0] wire_1;
  wire [0:0] wire_2;
  wire [7:0] wire_3;
  wire [0:0] wire_4;
  wire [63:0] wire_5;
  wire [63:0] wire_6;
  wire [0:0] wire_7;
  wire [7:0] wire_8;
  wire [0:0] wire_9;
  wire [63:0] wire_10;
  wire [0:0] wire_11;
  wire [7:0] wire_12;
  wire [63:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  wire [0:0] wire_16;
  wire [0:0] wire_17;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  wire [7:0] wire_20;
  wire [0:0] wire_21;
  wire [7:0] wire_22;
  wire [0:0] wire_23;
  wire [7:0] wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [7:0] wire_27;
  wire [7:0] wire_28;
  wire [0:0] wire_29;
  wire [7:0] wire_30;
  wire [7:0] wire_31;
  wire [0:0] wire_32;
  wire [7:0] wire_33;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  wire [7:0] wire_36;
  wire [0:0] wire_37;
  wire [7:0] wire_38;
  wire [7:0] wire_39;
  wire [0:0] wire_40;
  wire [0:0] wire_41;
  wire [0:0] wire_42;
  wire [0:0] wire_43;
  wire [0:0] wire_44;
  wire [0:0] wire_45;
  wire [63:0] wire_46;
  wire [0:0] wire_47;
  wire [0:0] wire_48;
  wire [0:0] wire_49;
  wire [0:0] wire_50;
  wire [0:0] wire_51;
  wire [0:0] wire_52;
  wire [0:0] wire_53;
  wire [0:0] wire_54;
  wire [0:0] wire_55;
  wire [0:0] wire_56;
  wire [0:0] wire_57;
  assign arch_input_enable = wire_57;
  wire [7:0] wire_58;
  wire [0:0] wire_59;
  wire [0:0] wire_60;
  wire [0:0] wire_61;
  wire [0:0] wire_62;
  wire [0:0] wire_63;
  wire [0:0] wire_64;
  wire [0:0] wire_65;
  wire [7:0] wire_66;
  wire [0:0] wire_67;
  wire [7:0] wire_68;
  wire [7:0] wire_69;
  wire [7:0] wire_70;
  wire [7:0] wire_71;
  wire [0:0] wire_72;
  wire [7:0] wire_73;
  wire [7:0] wire_74;
  wire [0:0] wire_75;
  wire [7:0] wire_76;
  wire [0:0] wire_77;
  wire [0:0] wire_78;
  wire [0:0] wire_79;
  wire [0:0] wire_80;
  wire [7:0] wire_81;
  wire [0:0] wire_82;
  wire [0:0] wire_83;
  wire [0:0] wire_84;
  wire [7:0] wire_85;
  wire [0:0] wire_86;
  wire [0:0] wire_87;
  assign arch_output_enable = wire_87;
  wire [0:0] wire_88;
  wire [0:0] wire_89;
  wire [0:0] wire_90;
  wire [7:0] wire_91;

endmodule
