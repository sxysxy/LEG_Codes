module _4zm16DatazmMUXzm8b (clk, rst, \�_____ , A3, A2, A1, A0, D0, D1, D2, D3, D4, D5, D6, D7, D8, D9, DA, DB, DC, DD, DE, DF, Output);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [0:0] \�_____ ;
  input  wire [0:0] A3;
  input  wire [0:0] A2;
  input  wire [0:0] A1;
  input  wire [0:0] A0;
  input  wire [7:0] D0;
  input  wire [7:0] D1;
  input  wire [7:0] D2;
  input  wire [7:0] D3;
  input  wire [7:0] D4;
  input  wire [7:0] D5;
  input  wire [7:0] D6;
  input  wire [7:0] D7;
  input  wire [7:0] D8;
  input  wire [7:0] D9;
  input  wire [7:0] DA;
  input  wire [7:0] DB;
  input  wire [7:0] DC;
  input  wire [7:0] DD;
  input  wire [7:0] DE;
  input  wire [7:0] DF;
  output  wire [7:0] Output;

  TC_Switch # (.UUID(64'd3168126685124603009 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_0 (.en(wire_15), .in(wire_27), .out(wire_1_11));
  TC_Switch # (.UUID(64'd2714236437993793899 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_1 (.en(wire_33), .in(wire_21), .out(wire_1_14));
  TC_Switch # (.UUID(64'd2115333001465120336 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_2 (.en(wire_34), .in(wire_22), .out(wire_1_5));
  TC_Switch # (.UUID(64'd972902543657377594 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_3 (.en(wire_12), .in(wire_37), .out(wire_1_13));
  TC_Switch # (.UUID(64'd3954311698125758584 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_4 (.en(wire_26), .in(wire_0), .out(wire_1_9));
  TC_Switch # (.UUID(64'd3029051993255470115 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_5 (.en(wire_24), .in(wire_4), .out(wire_1_2));
  TC_Switch # (.UUID(64'd935797790757251738 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_6 (.en(wire_13), .in(wire_10), .out(wire_1_1));
  TC_Switch # (.UUID(64'd2788006440996072909 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_7 (.en(wire_19), .in(wire_2), .out(wire_1_4));
  TC_Switch # (.UUID(64'd3349302701920232630 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_8 (.en(wire_9), .in(wire_18), .out(wire_1_3));
  TC_Switch # (.UUID(64'd1474541766342603399 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_9 (.en(wire_20), .in(wire_23), .out(wire_1_15));
  TC_Switch # (.UUID(64'd3566644400086355253 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_10 (.en(wire_6), .in(wire_16), .out(wire_1_10));
  TC_Switch # (.UUID(64'd998062770594250407 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_11 (.en(wire_31), .in(wire_11), .out(wire_1_0));
  TC_Switch # (.UUID(64'd4543826470152472504 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_12 (.en(wire_3), .in(wire_7), .out(wire_1_7));
  TC_Switch # (.UUID(64'd1165673664591012872 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_13 (.en(wire_17), .in(wire_8), .out(wire_1_8));
  TC_Switch # (.UUID(64'd2894624507190072279 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_14 (.en(wire_5), .in(wire_36), .out(wire_1_12));
  TC_Switch # (.UUID(64'd802842499667235992 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_15 (.en(wire_32), .in(wire_30), .out(wire_1_6));
  TC_Constant # (.UUID(64'd3308725179153905330 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_16 (.out());
  TC_Constant # (.UUID(64'd1816611684463819271 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_17 (.out());
  TC_Constant # (.UUID(64'd2843098605387643101 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_18 (.out());
  TC_Constant # (.UUID(64'd637348702270822651 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_19 (.out());
  TC_Constant # (.UUID(64'd203679650209229036 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_20 (.out());
  TC_Constant # (.UUID(64'd757784161449603171 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_21 (.out());
  TC_Constant # (.UUID(64'd775495168227954981 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_22 (.out());
  TC_Constant # (.UUID(64'd1543927474542086864 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_23 (.out());
  TC_Constant # (.UUID(64'd4031929066983585913 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_24 (.out());
  TC_Constant # (.UUID(64'd1895916469102550197 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_25 (.out());
  TC_Constant # (.UUID(64'd2523222794437694002 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_26 (.out());
  TC_Constant # (.UUID(64'd4004434000865767068 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_27 (.out());
  TC_Constant # (.UUID(64'd2023922848258811707 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_28 (.out());
  TC_Constant # (.UUID(64'd612582011967941220 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_29 (.out());
  _4zm16Selector # (.UUID(64'd3049110683819268068 ^ UUID)) _4zm16Selector_30 (.clk(clk), .rst(rst), .\�_____ (wire_25), .A3(wire_28), .A2(wire_29), .A1(wire_35), .A0(wire_14), .\0 (wire_15), .\1 (wire_33), .\2 (wire_34), .\3 (wire_12), .\4 (wire_26), .\5 (wire_24), .\6 (wire_13), .\7 (wire_19), .\8 (wire_32), .\9 (wire_5), .A(wire_17), .B(wire_3), .C(wire_31), .D(wire_6), .E(wire_20), .F(wire_9));

  wire [7:0] wire_0;
  assign wire_0 = D4;
  wire [7:0] wire_1;
  wire [7:0] wire_1_0;
  wire [7:0] wire_1_1;
  wire [7:0] wire_1_2;
  wire [7:0] wire_1_3;
  wire [7:0] wire_1_4;
  wire [7:0] wire_1_5;
  wire [7:0] wire_1_6;
  wire [7:0] wire_1_7;
  wire [7:0] wire_1_8;
  wire [7:0] wire_1_9;
  wire [7:0] wire_1_10;
  wire [7:0] wire_1_11;
  wire [7:0] wire_1_12;
  wire [7:0] wire_1_13;
  wire [7:0] wire_1_14;
  wire [7:0] wire_1_15;
  assign wire_1 = wire_1_0|wire_1_1|wire_1_2|wire_1_3|wire_1_4|wire_1_5|wire_1_6|wire_1_7|wire_1_8|wire_1_9|wire_1_10|wire_1_11|wire_1_12|wire_1_13|wire_1_14|wire_1_15;
  assign Output = wire_1;
  wire [7:0] wire_2;
  assign wire_2 = D7;
  wire [0:0] wire_3;
  wire [7:0] wire_4;
  assign wire_4 = D5;
  wire [0:0] wire_5;
  wire [0:0] wire_6;
  wire [7:0] wire_7;
  assign wire_7 = DB;
  wire [7:0] wire_8;
  assign wire_8 = DA;
  wire [0:0] wire_9;
  wire [7:0] wire_10;
  assign wire_10 = D6;
  wire [7:0] wire_11;
  assign wire_11 = DC;
  wire [0:0] wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  assign wire_14 = A0;
  wire [0:0] wire_15;
  wire [7:0] wire_16;
  assign wire_16 = DD;
  wire [0:0] wire_17;
  wire [7:0] wire_18;
  assign wire_18 = DF;
  wire [0:0] wire_19;
  wire [0:0] wire_20;
  wire [7:0] wire_21;
  assign wire_21 = D1;
  wire [7:0] wire_22;
  assign wire_22 = D2;
  wire [7:0] wire_23;
  assign wire_23 = DE;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  assign wire_25 = \�_____ ;
  wire [0:0] wire_26;
  wire [7:0] wire_27;
  assign wire_27 = D0;
  wire [0:0] wire_28;
  assign wire_28 = A3;
  wire [0:0] wire_29;
  assign wire_29 = A2;
  wire [7:0] wire_30;
  assign wire_30 = D8;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  assign wire_35 = A1;
  wire [7:0] wire_36;
  assign wire_36 = D9;
  wire [7:0] wire_37;
  assign wire_37 = D3;

endmodule
