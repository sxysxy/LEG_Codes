module RegisterFiles4x4zm8bzmEX (clk, rst, R_ADDR2, R_ADDR1, \input , W, W_ADDR, READ_2, READ_1);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [7:0] R_ADDR2;
  input  wire [7:0] R_ADDR1;
  input  wire [7:0] \input ;
  input  wire [0:0] W;
  input  wire [7:0] W_ADDR;
  output  wire [7:0] READ_2;
  output  wire [7:0] READ_1;

  TC_Splitter8 # (.UUID(64'd882782745428152396 ^ UUID)) Splitter8_0 (.in(wire_2), .out0(wire_31), .out1(wire_19), .out2(wire_41), .out3(wire_43), .out4(), .out5(), .out6(), .out7());
  TC_Not # (.UUID(64'd2853713365917981239 ^ UUID), .BIT_WIDTH(64'd1)) Not_1 (.in(wire_51), .out(wire_21));
  TC_Not # (.UUID(64'd1261395480174859567 ^ UUID), .BIT_WIDTH(64'd1)) Not_2 (.in(1'd0), .out());
  TC_Splitter8 # (.UUID(64'd1973127687343555926 ^ UUID)) Splitter8_3 (.in(wire_12), .out0(wire_35), .out1(wire_29), .out2(wire_34), .out3(wire_23), .out4(), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd3079115794087519115 ^ UUID)) Splitter8_4 (.in(wire_48), .out0(wire_49), .out1(wire_33), .out2(wire_52), .out3(wire_45), .out4(), .out5(), .out6(), .out7());
  TC_Constant # (.UUID(64'd1337279156297376405 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_5 (.out());
  TC_Constant # (.UUID(64'd1504053604124100900 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_6 (.out());
  TC_Constant # (.UUID(64'd197185958993143421 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_7 (.out());
  TC_Constant # (.UUID(64'd1305077583122413665 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_8 (.out());
  TC_Constant # (.UUID(64'd262881175941445387 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_9 (.out());
  TC_Constant # (.UUID(64'd2379093974745084274 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_10 (.out());
  TC_Constant # (.UUID(64'd1222797833592236955 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_11 (.out());
  TC_Constant # (.UUID(64'd2603573725252172514 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_12 (.out());
  TC_Constant # (.UUID(64'd2888588006610617179 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_13 (.out());
  TC_Constant # (.UUID(64'd1478113334755716975 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_14 (.out());
  TC_Constant # (.UUID(64'd835131139853149211 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_15 (.out());
  TC_Constant # (.UUID(64'd1688177124371010980 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_16 (.out());
  TC_Constant # (.UUID(64'd3613330890452583506 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_17 (.out());
  TC_Constant # (.UUID(64'd3302628028046420806 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_18 (.out());
  TC_Constant # (.UUID(64'd4249269848833075521 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_19 (.out());
  TC_Constant # (.UUID(64'd3596508173963038172 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_20 (.out());
  TC_Constant # (.UUID(64'd2717488093640686367 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_21 (.out());
  TC_Constant # (.UUID(64'd2102331319310393840 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_22 (.out());
  TC_Constant # (.UUID(64'd2687081266769874062 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_23 (.out());
  TC_Constant # (.UUID(64'd1606586793223473140 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_24 (.out());
  TC_Constant # (.UUID(64'd2252674971382543483 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_25 (.out());
  TC_Constant # (.UUID(64'd2306417731205294501 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_26 (.out());
  TC_Constant # (.UUID(64'd98213262110029667 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_27 (.out());
  TC_Constant # (.UUID(64'd4579190319189674387 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_28 (.out());
  RegisterPlus # (.UUID(64'd4411170466903339909 ^ UUID)) RegisterPlus_29 (.clk(clk), .rst(rst), .\�_____ (1'd0), .\�___________ (wire_6), .\�_____ (wire_42), .\�___________ (wire_0), .Output());
  RegisterPlus # (.UUID(64'd1518454392341965663 ^ UUID)) RegisterPlus_30 (.clk(clk), .rst(rst), .\�_____ (1'd0), .\�___________ (wire_6), .\�_____ (wire_47), .\�___________ (wire_15), .Output());
  RegisterPlus # (.UUID(64'd2141083928128949461 ^ UUID)) RegisterPlus_31 (.clk(clk), .rst(rst), .\�_____ (1'd0), .\�___________ (wire_6), .\�_____ (wire_16), .\�___________ (wire_17), .Output());
  RegisterPlus # (.UUID(64'd2927393123504819294 ^ UUID)) RegisterPlus_32 (.clk(clk), .rst(rst), .\�_____ (1'd0), .\�___________ (wire_6), .\�_____ (wire_4), .\�___________ (wire_22), .Output());
  RegisterPlus # (.UUID(64'd1096463846567443412 ^ UUID)) RegisterPlus_33 (.clk(clk), .rst(rst), .\�_____ (1'd0), .\�___________ (wire_6), .\�_____ (wire_24), .\�___________ (wire_5), .Output(wire_10));
  RegisterPlus # (.UUID(64'd3230815698680122166 ^ UUID)) RegisterPlus_34 (.clk(clk), .rst(rst), .\�_____ (1'd0), .\�___________ (wire_6), .\�_____ (wire_20), .\�___________ (wire_30), .Output());
  RegisterPlus # (.UUID(64'd2850840635606122746 ^ UUID)) RegisterPlus_35 (.clk(clk), .rst(rst), .\�_____ (1'd0), .\�___________ (wire_6), .\�_____ (wire_28), .\�___________ (wire_37), .Output());
  RegisterPlus # (.UUID(64'd23129690446293640 ^ UUID)) RegisterPlus_36 (.clk(clk), .rst(rst), .\�_____ (1'd0), .\�___________ (wire_6), .\�_____ (wire_11), .\�___________ (wire_13), .Output());
  RegisterPlus # (.UUID(64'd3555277572096861433 ^ UUID)) RegisterPlus_37 (.clk(clk), .rst(rst), .\�_____ (1'd0), .\�___________ (wire_6), .\�_____ (wire_39), .\�___________ (wire_9), .Output());
  RegisterPlus # (.UUID(64'd3280081926758671752 ^ UUID)) RegisterPlus_38 (.clk(clk), .rst(rst), .\�_____ (1'd0), .\�___________ (wire_6), .\�_____ (wire_44), .\�___________ (wire_7), .Output());
  RegisterPlus # (.UUID(64'd1796102896709818003 ^ UUID)) RegisterPlus_39 (.clk(clk), .rst(rst), .\�_____ (1'd0), .\�___________ (wire_6), .\�_____ (wire_32), .\�___________ (wire_1), .Output());
  RegisterPlus # (.UUID(64'd2486687895541499294 ^ UUID)) RegisterPlus_40 (.clk(clk), .rst(rst), .\�_____ (1'd0), .\�___________ (wire_6), .\�_____ (wire_40), .\�___________ (wire_46), .Output());
  RegisterPlus # (.UUID(64'd3757483585665027423 ^ UUID)) RegisterPlus_41 (.clk(clk), .rst(rst), .\�_____ (1'd0), .\�___________ (wire_6), .\�_____ (wire_26), .\�___________ (wire_3), .Output());
  RegisterPlus # (.UUID(64'd4538933183306051984 ^ UUID)) RegisterPlus_42 (.clk(clk), .rst(rst), .\�_____ (1'd0), .\�___________ (wire_6), .\�_____ (wire_27), .\�___________ (wire_25), .Output());
  RegisterPlus # (.UUID(64'd4077965182025163289 ^ UUID)) RegisterPlus_43 (.clk(clk), .rst(rst), .\�_____ (1'd0), .\�___________ (wire_6), .\�_____ (wire_36), .\�___________ (wire_18), .Output());
  _4zm16Selector # (.UUID(64'd527462030932968719 ^ UUID)) _4zm16Selector_44 (.clk(clk), .rst(rst), .\�_____ (wire_21), .A3(wire_43), .A2(wire_41), .A1(wire_19), .A0(wire_31), .\0 (wire_40), .\1 (wire_36), .\2 (wire_26), .\3 (wire_27), .\4 (wire_11), .\5 (wire_39), .\6 (wire_44), .\7 (wire_32), .\8 (wire_42), .\9 (wire_47), .A(wire_16), .B(wire_4), .C(wire_24), .D(wire_20), .E(wire_28), .F(wire_14));
  _4zm16DatazmMUXzm8b # (.UUID(64'd4055267262461330249 ^ UUID)) _4zm16DatazmMUXzm8b_45 (.clk(clk), .rst(rst), .\�_____ (1'd0), .A3(wire_45), .A2(wire_52), .A1(wire_33), .A0(wire_49), .D0(wire_46), .D1(wire_18), .D2(wire_3), .D3(wire_25), .D4(wire_13), .D5(wire_9), .D6(wire_7), .D7(wire_1), .D8(wire_0), .D9(wire_15), .DA(wire_17), .DB(wire_22), .DC(wire_10), .DD(wire_30), .DE(wire_37), .DF({{7{1'b0}}, wire_8 }), .Output(wire_38));
  _4zm16DatazmMUXzm8b # (.UUID(64'd1174776228594855952 ^ UUID)) _4zm16DatazmMUXzm8b_46 (.clk(clk), .rst(rst), .\�_____ (1'd0), .A3(wire_23), .A2(wire_34), .A1(wire_29), .A0(wire_35), .D0(wire_46), .D1(wire_18), .D2(wire_3), .D3(wire_25), .D4(wire_13), .D5(wire_9), .D6(wire_7), .D7(wire_1), .D8(wire_0), .D9(wire_15), .DA(wire_17), .DB(wire_22), .DC(wire_5), .DD(wire_30), .DE(wire_37), .DF({{7{1'b0}}, wire_8 }), .Output(wire_50));
  TC_Constant # (.UUID(64'd3975288366337731559 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd0)) Off_47 (.out(wire_8));

  wire [7:0] wire_0;
  wire [7:0] wire_1;
  wire [7:0] wire_2;
  assign wire_2 = W_ADDR;
  wire [7:0] wire_3;
  wire [0:0] wire_4;
  wire [7:0] wire_5;
  wire [7:0] wire_6;
  assign wire_6 = \input ;
  wire [7:0] wire_7;
  wire [0:0] wire_8;
  wire [7:0] wire_9;
  wire [7:0] wire_10;
  wire [0:0] wire_11;
  wire [7:0] wire_12;
  assign wire_12 = R_ADDR2;
  wire [7:0] wire_13;
  wire [0:0] wire_14;
  wire [7:0] wire_15;
  wire [0:0] wire_16;
  wire [7:0] wire_17;
  wire [7:0] wire_18;
  wire [0:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [7:0] wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [7:0] wire_25;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  wire [7:0] wire_30;
  wire [0:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  wire [0:0] wire_36;
  wire [7:0] wire_37;
  wire [7:0] wire_38;
  assign READ_1 = wire_38;
  wire [0:0] wire_39;
  wire [0:0] wire_40;
  wire [0:0] wire_41;
  wire [0:0] wire_42;
  wire [0:0] wire_43;
  wire [0:0] wire_44;
  wire [0:0] wire_45;
  wire [7:0] wire_46;
  wire [0:0] wire_47;
  wire [7:0] wire_48;
  assign wire_48 = R_ADDR1;
  wire [0:0] wire_49;
  wire [7:0] wire_50;
  assign READ_2 = wire_50;
  wire [0:0] wire_51;
  assign wire_51 = W;
  wire [0:0] wire_52;

endmodule
